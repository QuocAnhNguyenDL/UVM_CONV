`ifndef CONV_DEFINES
`define CONV_DEFINES


  `define COL 5
  `define BIT_WIDTH 8
  `define IN_WIDTH 8
  `define OUT_WIDTH 32
  `define IMG_SIZE 32

`endif